xph2sei412@cimeld18.4332:1491565437