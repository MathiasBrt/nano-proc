xph2sei412@cimeld20.4185:1492171606